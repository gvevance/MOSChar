NMOS characterisation

*************************************
* Include model file 
*************************************
.include 130nm_bulk.pm

*************************************
* Defining arameters 
*************************************
.param len = 0.3u
.param width = 100u 
.param lmin = 0.13u

*************************************
* Circuit definition
*************************************
vdd 1 0 dc 1.3
i0 2 1 dc 100
vds_ref 4 0 dc 0.2
e_amp 3 0 2 4 1e4
M1 2 3 0 0 nmos l={len} w={width} as={2*lmin*width} ad={2*lmin*width} ps={4*lmin+2*width} pd={4*lmin+2*width}


*************************************
* Control section
*************************************

.control 

save @M1[vdsat], @M1[vth], @M1[cgs], @M1[cgg],
+ @M1[gm], @M1[gds], @M1[gmbs], @M1[vsat]

* parameter sweep of width

let wmin = 10u
let wmax = 100u
let delta_w = 5u
let w = wmin

set filetype=ascii
set wr_singlescale
*set wr_vecnames

* loop
while w le wmax
    alter width w
    op
    wrdata values_nmos_v2_b.txt w, @M1[vdsat], @M1[cgs], @M1[cgg] 
    + @M1[gm], @M1[gds], @M1[gmbs], @M1[vth], @M1[vgs]
    set appendwrite
    let w = w + delta_w
end

* Run the sim
run

*wrdata values_nmos_v2_b.txt @M1[vdsat], @M1[cgs], @M1[cgg] 
*+ @M1[gm], @M1[gds], @M1[gmbs], @M1[vth], @M1[vgs]

* Plot commands
* plot @M1[id]
* plot @M1[gm]
* plot @M1[gmbs]
* plot @M1[gds]
* plot @M1[cgs]
* plot @M1[cgg]
* plot @M1[vdsat]
* plot @M1[vsat]


exit
.endc

*************************************
* End of file
*************************************
.end
