NMOS characterisation

*************************************
* Include model file 
*************************************
.include /home/gabriel/Desktop/Git/MOSChar/Model_files/130nm_bulk.pm

*************************************
* Defining arameters 
*************************************
.param len = 1.04u
.param width = 100u 
.param lmin = 0.13u

*************************************
* Circuit definition
*************************************
vdd 1 0 dc 1.3
i0 1 2 dc 100u
vds_ref 4 0 dc 0.2
e_amp 3 0 2 4 1e4
M1 2 3 0 0 nmos l={len} w={width} as={2*lmin*width} ad={2*lmin*width} ps={4*lmin+2*width} pd={4*lmin+2*width}


*************************************
* Control section
*************************************

.control 

* parameter sweep of width

let wmin = 30u
let wmax = 700u
let delta_w = 5u
let w = wmin

set filetype=ascii

save @M1[vdsat], @M1[vth], @M1[cgs], @M1[cgg],
+ @M1[gm], @M1[gds], @M1[gmbs], @M1[vsat]

echo "@M1[w] @M1[vgs] @M1[gm] @M1[gds] @M1[vdsat] @M1[vth] @M1[cgs] @M1[cgg] @M1[gmbs]" > /home/gabriel/Desktop/Git/MOSChar/tmp/values_nmos_v2_b.txt

* loop
while w le wmax
    
    * alter changes device value or device property ( not variables )
    alter @m1[w] = w
    
    * specify type of analysis
    op
    
    let gm = @M1[gm]
    let gds = @M1[gds]
    let vdsat = @M1[vdsat]
    let vgs = @M1[vgs]
    let vth = @M1[vth]
    let cgs = @M1[cgs]
    let cgg = @M1[cgg]
    let gmbs = @M1[gmbs]

    * run the sim
    run

    * append (>>) to file 
    echo "$&w" "$&vgs" "$&gm" "$&gds" "$&vdsat" "$&vth" "$&cgs" "$&cgg" "$&gmbs">> /home/gabriel/Desktop/Git/MOSChar/tmp/values_nmos_v2_b.txt
    
    * update variable w
    let w = w + delta_w

end

exit
.endc

*************************************
* End of file
*************************************
.end
