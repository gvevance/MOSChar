NMOS gm/ID circuit

.include 130nm_bulk.pm

* Parameters 
.param len=0.13u width=1.3u lmin=0.13u

* Circuit definition
vgs 1 0 dc 1
vds 2 0 dc 1
mn 2 1 0 0 NMOS l={len} w={width} ad={2*lmin*width} as={2*lmin*width} ps={4*lmin+1*width} pd={4*lmin+1*width}

.dc vgs 0 1.3 0.001

.control 

run

plot @mn[igs] @mn[id]

.endc
.end